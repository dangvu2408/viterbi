module ham_d (clk, rst, en_brch, data, hamd_1, hamd_2, hamd_3, hamd_4, hamd_5, hamd_6, hamd_7, hamd_8);

endmodule